/* alu
 * By: John Jekel
 *
 * ALU for the cpu
 *
*/

//TODO
