package common;
    typedef enum logic [7:0] {RASTER_CMD_NOP, RASTER_CMD_FILL, RASTER_CMD_POINT, RASTER_CMD_LINE /* TODO add others */} raster_command_t;
endpackage
