/* agu
 * By: John Jekel
 *
 * AGU for the cpu
 *
*/

module agu (

);

endmodule
