/* sp
 * By: John Jekel
 *
 * Stack pointer and the SP ALU for the cpu
 *
*/

//TODO
