/* rasterizer_controller
 * By: John Jekel
 *
 * CPU module for communicating the the rasterizer
 *
*/

module rasterizer_controller
    //import common::raster_command_t;
(
    /*
    input raster_command_t gpu_command,
    input logic [7:0] r4, r5, r6, r7,
    input logic [7:0] immediate,
    input logic gpu_submit,
    output logic gpu_busy,

    //CPU-GPU Interface
    rasterizer_if.cpu gpu_if
    */
);

//TODO

endmodule
