/* rasterizer_controller
 * By: John Jekel
 *
 * CPU module for communicating the the rasterizer
 *
*/

module rasterizer_controller
    import common::raster_command_t;
(

    //CPU-GPU Interface
    rasterizer_if.cpu gpu_if,
);

//TODO

endmodule
