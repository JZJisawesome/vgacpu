package common;
    typedef enum logic [7:0] {RASTER_CMD_NOP, RASTER_CMD_FILL, RASTER_CMD_POINT /* TODO add others */} raster_command_t;//TODO move this to some common package
endpackage
