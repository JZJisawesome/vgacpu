/* snd_controller
 * By: John Jekel
 *
 * CPU module for communicating the the sound module
 *
*/

module snd_controller (

);

//TODO

endmodule
