/* rasterizer_controller
 * By: John Jekel
 *
 * CPU module for communicating the the rasterizer
 *
*/

module rasterizer_controller (

);

//TODO

endmodule
