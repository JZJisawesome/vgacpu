/* vga
 * By: John Jekel
 *
 * Module for outputing VGA video from a framebuffer.
 *
*/
module vga
(
    input logic clk,//50MHz
    input logic n_rst,

    //VGA Outputs (640x480)
    output logic vga_r, vga_g, vga_b,
    output logic vga_hsync, vga_vsync

    //Framebuffer access
    //TODO
);

//TODO

endmodule
