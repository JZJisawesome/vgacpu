/* rf_mux
 * By: John Jekel
 *
 * Input multiplexer for the register file
 *
*/

//TODO
