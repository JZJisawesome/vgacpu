/* vgacpu
 * By: John Jekel
 *
 * Main module for the CPU in the hardware.
 *
*/
