/* pr
 * By: John Jekel
 *
 * Page register for the CPU
 *
*/

module pr (
    //TODO
);

endmodule
