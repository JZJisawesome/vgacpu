/* decode
 * By: John Jekel
 *
 * Decode unit for the cpu
 *
*/

//TODO
