/* sp
 * By: John Jekel
 *
 * Stack pointer and the SP ALU for the cpu
 *
*/

module sp (
    input clk,

    //TODO control signals: increment, decrement, stay the same, etc

    output [13:0] sp_addr

);

endmodule
