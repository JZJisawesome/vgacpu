/* fetch
 * By: John Jekel
 *
 * Fetch unit for the CPU
 *
*/

//TODO
