/* rf_mux
 * By: John Jekel
 *
 * Input multiplexer for the register file
 *
*/

module rf_mux (

    //TODO inputs

    output [7:0] rf_in

);

endmodule
