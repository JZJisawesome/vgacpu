/* fetch
 * By: John Jekel
 *
 * Fetch unit for the CPU
 *
*/

module fetch (
    input clk,
    input rst_async

);

endmodule
