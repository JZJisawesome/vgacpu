/* agu
 * By: John Jekel
 *
 * AGU for the cpu
 *
*/

//TODO
