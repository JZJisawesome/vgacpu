/* buttons_controller
 * By: John Jekel
 *
 * CPU module for reading the buttons
 *
*/

module button_controller (

);

//TODO

endmodule
