/* reg_file
 * By: John Jekel
 *
 * Register file for the CPU
 *
*/

module reg_file (
    input logic clk,

    //TODO control lines

    input logic [7:0] r_in,
    output logic [7:0] r0,
    output logic [7:0] r1,
    output logic [7:0] r4,
    output logic [7:0] r5,
    output logic [7:0] r6,
    output logic [7:0] r7,
    output logic [7:0] rX
);

//TODO

endmodule
